.PS
cct_init
ifdef(`NAND_gate',,`include(HOMELIB_`'liblog.m4)')
log_init

dim = 0.75

define( `mirror',`[
  line right_ dim*6/3
  "$V_{GS} = V_{DSsat} - V_{TH}$" at last line.c above
  M2: c_fet( up_ dim,,,) with .G at last line.end; rlabel( , "$M_2$");
  M4: c_fet( up_ dim,,,) with .S at M2.D; rlabel( , "$M_4$")
  line from M4.G left_ dim*6/3
  "$V_{G4} = 2V_{DSsat} + V_{TH}$" at last line.c above

  ground(at M2.S)
  arrow <- from M2.D right dim/2 up dim/6
  "$V_{DSsat}$" above ljust

  arrow <- from M4.D right dim/2 up dim/6
  "$\geq 2 V_{DSsat}$" above ljust

  line from M4.D up_ dim/4
]')

M: mirror

.PE